// This is a wrapper for the SimdPermutation module
module SimdPermWrapper import rvv_pkg::*; #(
    parameter int NumLanes = 8,
    parameter int NumSegments = 8,
    parameter int NumRotationRadix = 4,
    parameter int SizeXbar = 32,
    // DO NOT CHANGE!
    parameter int XLEN = 64,
    parameter int NumBanks = 8,
    parameter int UsePipeline = 1,
    parameter int NumInOuts = NumLanes * NumBanks
) (
   // Declare some signals so we can see how I/O works
   input              clk_i,
   input              rst_ni,

   input              operand_valid_i,
   output             operand_ready_o,
   input              selIdxVal,
   input              [XLEN-1:0] [NumInOuts-1:0] operand_i,

   input              permute_i,
   input              vlut_e lut_mode_i,

   input              result_ready_i,
   output             result_valid_o,
   output             [XLEN-1:0] [NumInOuts-1:0] result_o 
);

   // dut
   SimdPermutation simd_permutation(
    .clock(clk_i),
    .reset(~rst_ni),

    .io_inValid(operand_valid_i),
    .io_inReady(operand_ready_o),
    .io_selIdxVal(selIdxVal),

    .io_inData_0_0(operand_i[0]),
    .io_inData_0_1(operand_i[1]),
    .io_inData_0_2(operand_i[2]),
    .io_inData_0_3(operand_i[3]),
    .io_inData_0_4(operand_i[4]),
    .io_inData_0_5(operand_i[5]),
    .io_inData_0_6(operand_i[6]),
    .io_inData_0_7(operand_i[7]),
    .io_inData_1_0(operand_i[8]),
    .io_inData_1_1(operand_i[9]),
    .io_inData_1_2(operand_i[10]),
    .io_inData_1_3(operand_i[11]),
    .io_inData_1_4(operand_i[12]),
    .io_inData_1_5(operand_i[13]),
    .io_inData_1_6(operand_i[14]),
    .io_inData_1_7(operand_i[15]),
    .io_inData_2_0(operand_i[16]),
    .io_inData_2_1(operand_i[17]),
    .io_inData_2_2(operand_i[18]),
    .io_inData_2_3(operand_i[19]),
    .io_inData_2_4(operand_i[20]),
    .io_inData_2_5(operand_i[21]),
    .io_inData_2_6(operand_i[22]),
    .io_inData_2_7(operand_i[23]),
    .io_inData_3_0(operand_i[24]),
    .io_inData_3_1(operand_i[25]),
    .io_inData_3_2(operand_i[26]),
    .io_inData_3_3(operand_i[27]),
    .io_inData_3_4(operand_i[28]),
    .io_inData_3_5(operand_i[29]),
    .io_inData_3_6(operand_i[30]),
    .io_inData_3_7(operand_i[31]),
    .io_inData_4_0(operand_i[32]),
    .io_inData_4_1(operand_i[33]),
    .io_inData_4_2(operand_i[34]),
    .io_inData_4_3(operand_i[35]),
    .io_inData_4_4(operand_i[36]),
    .io_inData_4_5(operand_i[37]),
    .io_inData_4_6(operand_i[38]),
    .io_inData_4_7(operand_i[39]),
    .io_inData_5_0(operand_i[40]),
    .io_inData_5_1(operand_i[41]),
    .io_inData_5_2(operand_i[42]),
    .io_inData_5_3(operand_i[43]),
    .io_inData_5_4(operand_i[44]),
    .io_inData_5_5(operand_i[45]),
    .io_inData_5_6(operand_i[46]),
    .io_inData_5_7(operand_i[47]),
    .io_inData_6_0(operand_i[48]),
    .io_inData_6_1(operand_i[49]),
    .io_inData_6_2(operand_i[50]),
    .io_inData_6_3(operand_i[51]),
    .io_inData_6_4(operand_i[52]),
    .io_inData_6_5(operand_i[53]),
    .io_inData_6_6(operand_i[54]),
    .io_inData_6_7(operand_i[55]),
    .io_inData_7_0(operand_i[56]),
    .io_inData_7_1(operand_i[57]),
    .io_inData_7_2(operand_i[58]),
    .io_inData_7_3(operand_i[59]),
    .io_inData_7_4(operand_i[60]),
    .io_inData_7_5(operand_i[61]),
    .io_inData_7_6(operand_i[62]),
    .io_inData_7_7(operand_i[63]),

    .io_permute(permute_i),
    .io_mode(lut_mode_i), 
    .io_outValid(result_valid_o), 
    .io_outReady(result_ready_i), 

    .io_outData_0_0(result_o[0]),
    .io_outData_0_1(result_o[1]),
    .io_outData_0_2(result_o[2]),
    .io_outData_0_3(result_o[3]),
    .io_outData_0_4(result_o[4]),
    .io_outData_0_5(result_o[5]),
    .io_outData_0_6(result_o[6]),
    .io_outData_0_7(result_o[7]),
    .io_outData_1_0(result_o[8]),
    .io_outData_1_1(result_o[9]),
    .io_outData_1_2(result_o[10]),
    .io_outData_1_3(result_o[11]),
    .io_outData_1_4(result_o[12]),
    .io_outData_1_5(result_o[13]),
    .io_outData_1_6(result_o[14]),
    .io_outData_1_7(result_o[15]),
    .io_outData_2_0(result_o[16]),
    .io_outData_2_1(result_o[17]),
    .io_outData_2_2(result_o[18]),
    .io_outData_2_3(result_o[19]),
    .io_outData_2_4(result_o[20]),
    .io_outData_2_5(result_o[21]),
    .io_outData_2_6(result_o[22]),
    .io_outData_2_7(result_o[23]),
    .io_outData_3_0(result_o[24]),
    .io_outData_3_1(result_o[25]),
    .io_outData_3_2(result_o[26]),
    .io_outData_3_3(result_o[27]),
    .io_outData_3_4(result_o[28]),
    .io_outData_3_5(result_o[29]),
    .io_outData_3_6(result_o[30]),
    .io_outData_3_7(result_o[31]),
    .io_outData_4_0(result_o[32]),
    .io_outData_4_1(result_o[33]),
    .io_outData_4_2(result_o[34]),
    .io_outData_4_3(result_o[35]),
    .io_outData_4_4(result_o[36]),
    .io_outData_4_5(result_o[37]),
    .io_outData_4_6(result_o[38]),
    .io_outData_4_7(result_o[39]),
    .io_outData_5_0(result_o[40]),
    .io_outData_5_1(result_o[41]),
    .io_outData_5_2(result_o[42]),
    .io_outData_5_3(result_o[43]),
    .io_outData_5_4(result_o[44]),
    .io_outData_5_5(result_o[45]),
    .io_outData_5_6(result_o[46]),
    .io_outData_5_7(result_o[47]),
    .io_outData_6_0(result_o[48]),
    .io_outData_6_1(result_o[49]),
    .io_outData_6_2(result_o[50]),
    .io_outData_6_3(result_o[51]),
    .io_outData_6_4(result_o[52]),
    .io_outData_6_5(result_o[53]),
    .io_outData_6_6(result_o[54]),
    .io_outData_6_7(result_o[55]),
    .io_outData_7_0(result_o[56]),
    .io_outData_7_1(result_o[57]),
    .io_outData_7_2(result_o[58]),
    .io_outData_7_3(result_o[59]),
    .io_outData_7_4(result_o[60]),
    .io_outData_7_5(result_o[61]),
    .io_outData_7_6(result_o[62]),
    .io_outData_7_7(result_o[63])
   );

endmodule

/home/whxu/code/chisel-simd-permutation/generated/SimdPermutation_2048_16.sv